 
	module bch_64_dec (
	clk,
	reset_n,
	enable,
	i_code,
	o_data,
	o_valid,
	o_err_corr,
	o_err_detec,
	o_err_fatal

	);

	//------ INPUT PORTS -----
	input clk ;
	input reset_n;
	input enable;
	input [0:77] i_code;


	//------OUTPUT PORTS -----
	output [0:63] o_data;
	output o_valid;
	output o_err_corr;
	output o_err_detec;
	output o_err_fatal;

	//---- INTERNAL VARIABLES ---

	reg [0:77] codereg ;
	reg o_err_fatal;
	reg o_err_detec;
	reg o_err_corr;
	reg o_valid;
	wire noerr; 
	wire [0:63] corr_word; 


	wire [0:13] synd ; 
	wire [0:63] flip ; // databits error mask 
	reg [0:63] o_data; 
	wire [0:63] data = codereg[14:77] ; //extract databits 
	

	//---STATEMENTS 
	 


	
//----------Syndrome Generation-------------//
assign synd[0] = codereg[0] ^ codereg[7] ^ codereg[11] ^ codereg[14] ^ codereg[15] ^ codereg[19] ^ codereg[21] ^ codereg[22] ^ codereg[23] ^ codereg[25] ^ codereg[27] ^ codereg[28] ^ codereg[30] ^ codereg[31] ^ codereg[37] ^ codereg[38] ^ codereg[41] ^ codereg[42] ^ codereg[44] ^ codereg[46] ^ codereg[49] ^ codereg[50] ^ codereg[51] ^ codereg[54] ^ codereg[55] ^ codereg[56] ^ codereg[57] ^ codereg[59] ^ codereg[60] ^ codereg[62] ^ codereg[67] ^ codereg[69] ^ codereg[71] ^ codereg[73] ^ codereg[74] ^ codereg[75] ^ codereg[76] ^ codereg[77];
assign synd[1] = codereg[1] ^ codereg[8] ^ codereg[12] ^ codereg[15] ^ codereg[16] ^ codereg[20] ^ codereg[22] ^ codereg[23] ^ codereg[24] ^ codereg[26] ^ codereg[28] ^ codereg[29] ^ codereg[31] ^ codereg[32] ^ codereg[38] ^ codereg[39] ^ codereg[42] ^ codereg[43] ^ codereg[45] ^ codereg[47] ^ codereg[50] ^ codereg[51] ^ codereg[52] ^ codereg[55] ^ codereg[56] ^ codereg[57] ^ codereg[58] ^ codereg[60] ^ codereg[61] ^ codereg[63] ^ codereg[68] ^ codereg[70] ^ codereg[72] ^ codereg[74] ^ codereg[75] ^ codereg[76] ^ codereg[77];
assign synd[2] = codereg[2] ^ codereg[9] ^ codereg[13] ^ codereg[16] ^ codereg[17] ^ codereg[21] ^ codereg[23] ^ codereg[24] ^ codereg[25] ^ codereg[27] ^ codereg[29] ^ codereg[30] ^ codereg[32] ^ codereg[33] ^ codereg[39] ^ codereg[40] ^ codereg[43] ^ codereg[44] ^ codereg[46] ^ codereg[48] ^ codereg[51] ^ codereg[52] ^ codereg[53] ^ codereg[56] ^ codereg[57] ^ codereg[58] ^ codereg[59] ^ codereg[61] ^ codereg[62] ^ codereg[64] ^ codereg[69] ^ codereg[71] ^ codereg[73] ^ codereg[75] ^ codereg[76] ^ codereg[77];
assign synd[3] = codereg[3] ^ codereg[7] ^ codereg[10] ^ codereg[11] ^ codereg[15] ^ codereg[17] ^ codereg[18] ^ codereg[19] ^ codereg[21] ^ codereg[23] ^ codereg[24] ^ codereg[26] ^ codereg[27] ^ codereg[33] ^ codereg[34] ^ codereg[37] ^ codereg[38] ^ codereg[40] ^ codereg[42] ^ codereg[45] ^ codereg[46] ^ codereg[47] ^ codereg[50] ^ codereg[51] ^ codereg[52] ^ codereg[53] ^ codereg[55] ^ codereg[56] ^ codereg[58] ^ codereg[63] ^ codereg[65] ^ codereg[67] ^ codereg[69] ^ codereg[70] ^ codereg[71] ^ codereg[72] ^ codereg[73] ^ codereg[75];
assign synd[4] = codereg[4] ^ codereg[8] ^ codereg[11] ^ codereg[12] ^ codereg[16] ^ codereg[18] ^ codereg[19] ^ codereg[20] ^ codereg[22] ^ codereg[24] ^ codereg[25] ^ codereg[27] ^ codereg[28] ^ codereg[34] ^ codereg[35] ^ codereg[38] ^ codereg[39] ^ codereg[41] ^ codereg[43] ^ codereg[46] ^ codereg[47] ^ codereg[48] ^ codereg[51] ^ codereg[52] ^ codereg[53] ^ codereg[54] ^ codereg[56] ^ codereg[57] ^ codereg[59] ^ codereg[64] ^ codereg[66] ^ codereg[68] ^ codereg[70] ^ codereg[71] ^ codereg[72] ^ codereg[73] ^ codereg[74] ^ codereg[76];
assign synd[5] = codereg[5] ^ codereg[9] ^ codereg[12] ^ codereg[13] ^ codereg[17] ^ codereg[19] ^ codereg[20] ^ codereg[21] ^ codereg[23] ^ codereg[25] ^ codereg[26] ^ codereg[28] ^ codereg[29] ^ codereg[35] ^ codereg[36] ^ codereg[39] ^ codereg[40] ^ codereg[42] ^ codereg[44] ^ codereg[47] ^ codereg[48] ^ codereg[49] ^ codereg[52] ^ codereg[53] ^ codereg[54] ^ codereg[55] ^ codereg[57] ^ codereg[58] ^ codereg[60] ^ codereg[65] ^ codereg[67] ^ codereg[69] ^ codereg[71] ^ codereg[72] ^ codereg[73] ^ codereg[74] ^ codereg[75] ^ codereg[77];
assign synd[6] = codereg[6] ^ codereg[10] ^ codereg[13] ^ codereg[14] ^ codereg[18] ^ codereg[20] ^ codereg[21] ^ codereg[22] ^ codereg[24] ^ codereg[26] ^ codereg[27] ^ codereg[29] ^ codereg[30] ^ codereg[36] ^ codereg[37] ^ codereg[40] ^ codereg[41] ^ codereg[43] ^ codereg[45] ^ codereg[48] ^ codereg[49] ^ codereg[50] ^ codereg[53] ^ codereg[54] ^ codereg[55] ^ codereg[56] ^ codereg[58] ^ codereg[59] ^ codereg[61] ^ codereg[66] ^ codereg[68] ^ codereg[70] ^ codereg[72] ^ codereg[73] ^ codereg[74] ^ codereg[75] ^ codereg[76];
assign synd[7] = codereg[0] ^ codereg[5] ^ codereg[7] ^ codereg[9] ^ codereg[10] ^ codereg[14] ^ codereg[17] ^ codereg[18] ^ codereg[19] ^ codereg[20] ^ codereg[23] ^ codereg[25] ^ codereg[28] ^ codereg[31] ^ codereg[33] ^ codereg[34] ^ codereg[36] ^ codereg[38] ^ codereg[40] ^ codereg[46] ^ codereg[47] ^ codereg[50] ^ codereg[55] ^ codereg[56] ^ codereg[57] ^ codereg[59] ^ codereg[61] ^ codereg[62] ^ codereg[63] ^ codereg[66] ^ codereg[67] ^ codereg[68] ^ codereg[72] ^ codereg[73] ^ codereg[75] ^ codereg[76];
assign synd[8] = codereg[4] ^ codereg[5] ^ codereg[8] ^ codereg[13] ^ codereg[14] ^ codereg[15] ^ codereg[17] ^ codereg[19] ^ codereg[20] ^ codereg[21] ^ codereg[24] ^ codereg[25] ^ codereg[26] ^ codereg[30] ^ codereg[31] ^ codereg[33] ^ codereg[34] ^ codereg[37] ^ codereg[38] ^ codereg[45] ^ codereg[49] ^ codereg[50] ^ codereg[51] ^ codereg[52] ^ codereg[53] ^ codereg[55] ^ codereg[58] ^ codereg[59] ^ codereg[61] ^ codereg[65] ^ codereg[67] ^ codereg[68] ^ codereg[69] ^ codereg[70] ^ codereg[72] ^ codereg[73] ^ codereg[75] ^ codereg[76] ^ codereg[77];
assign synd[9] = codereg[3] ^ codereg[7] ^ codereg[8] ^ codereg[9] ^ codereg[10] ^ codereg[11] ^ codereg[13] ^ codereg[16] ^ codereg[17] ^ codereg[19] ^ codereg[23] ^ codereg[25] ^ codereg[26] ^ codereg[27] ^ codereg[28] ^ codereg[30] ^ codereg[31] ^ codereg[33] ^ codereg[34] ^ codereg[35] ^ codereg[37] ^ codereg[38] ^ codereg[39] ^ codereg[40] ^ codereg[41] ^ codereg[42] ^ codereg[43] ^ codereg[48] ^ codereg[50] ^ codereg[52] ^ codereg[53] ^ codereg[57] ^ codereg[60] ^ codereg[61] ^ codereg[62] ^ codereg[63] ^ codereg[66] ^ codereg[68] ^ codereg[71] ^ codereg[74] ^ codereg[76] ^ codereg[77];
assign synd[10] = codereg[1] ^ codereg[5] ^ codereg[6] ^ codereg[7] ^ codereg[8] ^ codereg[9] ^ codereg[11] ^ codereg[14] ^ codereg[15] ^ codereg[17] ^ codereg[21] ^ codereg[23] ^ codereg[24] ^ codereg[25] ^ codereg[26] ^ codereg[28] ^ codereg[29] ^ codereg[31] ^ codereg[32] ^ codereg[33] ^ codereg[35] ^ codereg[36] ^ codereg[37] ^ codereg[38] ^ codereg[39] ^ codereg[40] ^ codereg[41] ^ codereg[46] ^ codereg[48] ^ codereg[50] ^ codereg[51] ^ codereg[55] ^ codereg[58] ^ codereg[59] ^ codereg[60] ^ codereg[61] ^ codereg[64] ^ codereg[66] ^ codereg[69] ^ codereg[72] ^ codereg[74] ^ codereg[75] ^ codereg[77];
assign synd[11] = codereg[4] ^ codereg[6] ^ codereg[8] ^ codereg[9] ^ codereg[13] ^ codereg[16] ^ codereg[17] ^ codereg[18] ^ codereg[19] ^ codereg[22] ^ codereg[24] ^ codereg[27] ^ codereg[30] ^ codereg[32] ^ codereg[33] ^ codereg[35] ^ codereg[37] ^ codereg[39] ^ codereg[45] ^ codereg[46] ^ codereg[49] ^ codereg[54] ^ codereg[55] ^ codereg[56] ^ codereg[58] ^ codereg[60] ^ codereg[61] ^ codereg[62] ^ codereg[65] ^ codereg[66] ^ codereg[67] ^ codereg[71] ^ codereg[72] ^ codereg[74] ^ codereg[75];
assign synd[12] = codereg[3] ^ codereg[4] ^ codereg[7] ^ codereg[12] ^ codereg[13] ^ codereg[14] ^ codereg[16] ^ codereg[18] ^ codereg[19] ^ codereg[20] ^ codereg[23] ^ codereg[24] ^ codereg[25] ^ codereg[29] ^ codereg[30] ^ codereg[32] ^ codereg[33] ^ codereg[36] ^ codereg[37] ^ codereg[44] ^ codereg[48] ^ codereg[49] ^ codereg[50] ^ codereg[51] ^ codereg[52] ^ codereg[54] ^ codereg[57] ^ codereg[58] ^ codereg[60] ^ codereg[64] ^ codereg[66] ^ codereg[67] ^ codereg[68] ^ codereg[69] ^ codereg[71] ^ codereg[72] ^ codereg[74] ^ codereg[75] ^ codereg[76];
assign synd[13] = codereg[2] ^ codereg[6] ^ codereg[7] ^ codereg[8] ^ codereg[9] ^ codereg[10] ^ codereg[12] ^ codereg[15] ^ codereg[16] ^ codereg[18] ^ codereg[22] ^ codereg[24] ^ codereg[25] ^ codereg[26] ^ codereg[27] ^ codereg[29] ^ codereg[30] ^ codereg[32] ^ codereg[33] ^ codereg[34] ^ codereg[36] ^ codereg[37] ^ codereg[38] ^ codereg[39] ^ codereg[40] ^ codereg[41] ^ codereg[42] ^ codereg[47] ^ codereg[49] ^ codereg[51] ^ codereg[52] ^ codereg[56] ^ codereg[59] ^ codereg[60] ^ codereg[61] ^ codereg[62] ^ codereg[65] ^ codereg[67] ^ codereg[70] ^ codereg[73] ^ codereg[75] ^ codereg[76];

wire ignore = (synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13]);

//----------Syndrome Decoding----------------//
assign noerr = ~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13];
assign flip[0] = (synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[1] = (synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[2] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[3] = (~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13]);
assign flip[4] = (~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[5] = (synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[6] = (~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[7] = (synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[8] = (synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[9] = (synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[10] = (~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[11] = (synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[12] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[13] = (synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[14] = (synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[15] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[16] = (synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[17] = (synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[18] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[19] = (~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[20] = (~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[21] = (~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13]);
assign flip[22] = (~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[23] = (synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[24] = (synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[25] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[26] = (~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[27] = (synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[28] = (synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[29] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[30] = (synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[31] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13]);
assign flip[32] = (synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13]);
assign flip[33] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[34] = (~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[35] = (synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[36] = (synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[37] = (synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[38] = (~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[39] = (~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[40] = (synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[41] = (synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13]);
assign flip[42] = (synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[43] = (synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[44] = (~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[45] = (synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[46] = (synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[47] = (~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[48] = (synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[49] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13]);
assign flip[50] = (~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[51] = (~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13]);
assign flip[52] = (~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[53] = (synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[54] = (~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[55] = (synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13]);
assign flip[56] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[57] = (synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[58] = (~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[59] = (synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13]);
assign flip[60] = (synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13]);
assign flip[61] = (synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13]);
assign flip[62] = (synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13]);
assign flip[63] = (synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13])|(synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & ~synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & ~synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & ~synd[10] & synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & ~synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & ~synd[4] & synd[5] & ~synd[6] & synd[7] & synd[8] & ~synd[9] & synd[10] & ~synd[11] & ~synd[12] & ~synd[13])|(synd[0] & synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & ~synd[6] & ~synd[7] & synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & ~synd[12] & synd[13])|(synd[0] & synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & synd[11] & synd[12] & synd[13])|(synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & ~synd[8] & synd[9] & ~synd[10] & ~synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & synd[5] & synd[6] & ~synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & ~synd[6] & ~synd[7] & synd[8] & ~synd[9] & synd[10] & synd[11] & synd[12] & ~synd[13])|(synd[0] & ~synd[1] & synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & synd[1] & ~synd[2] & synd[3] & synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & synd[10] & ~synd[11] & ~synd[12] & synd[13])|(~synd[0] & ~synd[1] & synd[2] & ~synd[3] & synd[4] & ~synd[5] & synd[6] & ~synd[7] & synd[8] & ~synd[9] & ~synd[10] & synd[11] & synd[12] & ~synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & synd[3] & ~synd[4] & ~synd[5] & synd[6] & synd[7] & ~synd[8] & synd[9] & ~synd[10] & synd[11] & synd[12] & synd[13])|(~synd[0] & ~synd[1] & ~synd[2] & ~synd[3] & synd[4] & synd[5] & synd[6] & synd[7] & ~synd[8] & ~synd[9] & synd[10] & ~synd[11] & synd[12] & synd[13]);



	

	assign corr_word = data[0:63] ^ flip[0:63]; 


	////////// REGISTER INPUT CODEWORD ////////////////

	always @(posedge clk or negedge reset_n) begin
		if (!reset_n) 
			// reset
			codereg <= 0 ;
		
		else if (enable)  
			codereg <= i_code; 
		 
	end

	//////////// GET OUTPUT ////////////////////////
	always @(posedge clk or negedge reset_n) begin
		if (!reset_n) begin
			// reset
			o_data <= 0;
			o_valid <= 0; 
			o_err_detec <=0;
			o_err_corr <= 0;
			o_err_fatal <= 0;
		end
		else if (enable) begin

			o_data <= corr_word ;
			o_err_detec <= ~noerr ;
			o_err_corr <= |flip ; // found one name match 
			o_err_fatal <= ~(|flip) & ~noerr & ~ignore; // has error AND syndrome has even parity. 2 err or more 
			o_valid <= 1 ; 
			
		end
	end



	endmodule 
	//--------- end of file ------//



	 
